--Rock Boynton
--Date: 10/30/17
--Course: CE 1901-021
--Professor: Dr. Livingston
--Purpose: This is the Structural VHDL for the Carry-Select Adder (CLA)
--         implementation adding two 8-bit numbers.

library IEEE;
use IEEE.std_logic_1164.all;