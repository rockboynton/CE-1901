----Rock Boynton
----Date: 10/30/17
----Course: CE 1901-021
----Professor: Dr. Livingston
----Purpose: This is the Full Adder component 
--
--library IEEE;
--use IEEE.std_logic_1164.all;
--
--entity CLA4 is 
--	port(Af: in std_logic;
--	     Bf: in std_logic;
--		  Cinf: in std_logic;
--		  Sf: out std_logic;
--		  Coutf: out std_logic);
--		  
--end entity CLA4;
--
--architecture SSTRUCTURAL of CLA4 is 
--
--signal G : std_logic_vector(3 downto 0);
--signal P : std_logic_vector(3 downto 0);
--
--begin
--
--
--
--end architecture DATAFLOW;
